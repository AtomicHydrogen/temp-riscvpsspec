package mulSat;
export  mulSat::*;
//USELESS FILE

    function Bit#(64) sixtSat (Bit#(64) rs1, Bit#(64) rs2);
        Bit#(64) outp;
        for (Integer i = 0; i < 4; i = i + 1);
            
        return outp;
    endfunction





endpackage